library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_misc.all;
  use IEEE.numeric_std.all;
  use work.roling_register_p.all;
  use work.xgen_axistream_32.all;
  use work.TX_DAC_control_pack.all;


entity TX_DAC_control_w_regInterface is
  generic ( 
    asicNumber : integer := 0
  );
  port (
    clk : std_logic;
    rst : std_logic;


    reg : registerT;


    TX_DAC_control_out : out  TX_DAC_control := TX_DAC_control_null
    
  );
end entity;

architecture rtl of TX_DAC_control_w_regInterface is

  
  
  
  signal  reg_data_m2s : axisStream_32_m2s := axisStream_32_m2s_null;  
  signal  reg_data_s2m : axisStream_32_s2m := axisStream_32_s2m_null;  





  signal   i_reg           :  registerT:= registerT_null;


begin

  DUT :  entity work.tx_dac_control_axi port map(
    clk => clk,
    regin => reg,
    reg_data_m2s => reg_data_m2s,
    reg_data_s2m => reg_data_s2m,
    sin  => TX_DAC_control_out.SIN,
    sclk => TX_DAC_control_out.SCLK,
    pclk => TX_DAC_control_out.PCLK
  );


  process(clk) is
    variable regTX : axisStream_32_master := axisStream_32_master_null;
    variable REG_DATA :  STD_LOGIC_VECTOR(31 downto 0) := (others => '0');
    variable TargetAsic : integer := 0;
  begin
    if rising_edge(clk) then 
      pull(regTx, reg_data_s2m);
			  TargetAsic :=  to_integer(unsigned(i_reg.address(15 downto 7)));
        if (TargetAsic = asicNumber + 1 or TargetAsic = 0)  and or_reduce(i_reg.address(6 downto 0)) = '1'  Then 
            REG_DATA := (others => '0');
            REG_DATA(18 downto 12) := std_logic_vector(unsigned( i_reg.address(6 downto 0)) - 1);
            REG_DATA(11 downto 0)  := i_reg.value(11 downto 0);
            send_data(regTX, REG_DATA);

        end if;
      push(regTx,reg_data_m2s);
    end if;
  end process;


  



  
  
  reg_buffer : entity work.registerBuffer generic map (
        Depth =>  10
  ) port map (
    
    clk =>clk,
    registersIn   => reg,
    registersOut  => i_reg
  );
end architecture;